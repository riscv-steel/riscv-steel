// ----------------------------------------------------------------------------
// Copyright (c) 2020-2024 RISC-V Steel contributors
//
// This work is licensed under the MIT License, see LICENSE file for details.
// SPDX-License-Identifier: MIT
// ----------------------------------------------------------------------------

module spi_cmod_a7 #( 

  parameter GPIO_WIDTH = 1,
  parameter SPI_NUM_CHIP_SELECT = 1

  )(

  input   wire clock,
  input   wire reset,
  input   wire uart_rx,
  output  wire uart_tx,
  output  wire sclk,
  output  wire pico,
  input   wire poci,
  output  wire cs

  );

  // Buttons debouncing
  reg reset_debounced;
  always @(posedge clock) begin
    reset_debounced <= reset;
  end

  rvsteel_mcu #(

    .CLOCK_FREQUENCY          (12000000               ),
    .UART_BAUD_RATE           (9600                   ),
    .MEMORY_SIZE              (131072                 ),
    .MEMORY_INIT_FILE         ("spi_demo.hex"         ),
    .BOOT_ADDRESS             (32'h00000000           ),
    .GPIO_WIDTH               (GPIO_WIDTH             ),
    .SPI_NUM_CHIP_SELECT      (SPI_NUM_CHIP_SELECT    )

  ) rvsteel_mcu_instance (

    .clock                    (clock                  ),
    .reset                    (reset_debounced        ),
    .halt                     (1'b0                   ),
    .uart_rx                  (uart_rx                ),
    .uart_tx                  (uart_tx                ),
    .gpio_input               ({GPIO_WIDTH{1'b0}}     ), // pull-down
    .gpio_oe                  (), // unused
    .gpio_output              (), // unused
    .sclk                     (sclk                   ),
    .pico                     (pico                   ),
    .poci                     (poci                   ),
    .cs                       (cs                     )

  );

endmodule