// ----------------------------------------------------------------------------
// Copyright (c) 2020-2024 RISC-V Steel contributors
//
// This work is licensed under the MIT License, see LICENSE file for details.
// SPDX-License-Identifier: MIT
// ----------------------------------------------------------------------------

module hello_world_cmod_a7 (

  input   wire clock,
  input   wire reset,
  output  wire uart_tx

  );

  // Push-button debouncing
  reg reset_debounced;
  always @(posedge clock) begin
    reset_debounced <= reset;
  end

  rvsteel_soc #(

  // Please adjust these two parameters accordingly

  .CLOCK_FREQUENCY          (12000000                   ),
  .MEMORY_INIT_FILE         ("hello_world.hex"          )

  ) rvsteel_soc_instance (

  // Note that unused inputs are hardwired to zero,
  // while unused outputs are left open.

  .clock                    (clock                      ),
  .reset                    (reset_debounced            ),
  .halt                     (1'b0                       ),
  .uart_rx                  (/* unused, leave open */   ),
  .uart_tx                  (uart_tx                    ),
  .gpio_input               (1'b0                       ),
  .gpio_oe                  (/* unused, leave open */   ),
  .gpio_output              (/* unused, leave open */   ),
  .sclk                     (/* unused, leave open */   ),
  .pico                     (/* unused, leave open */   ),
  .poci                     (1'b0                       ),
  .cs                       (/* unused, leave open */   )

  );

endmodule